// TCORE RISC-V Processor
// Copyright (c) 2024 Kerim TURAK
// Permission is hereby granted, free of charge, to any person obtaining a copy of this software
// and associated documentation files (the "Software"), to deal in the Software without restriction,
// including without limitation the rights to use, copy, modify, merge, publish, distribute,
// sublicense, and/or sell copies of the Software, and to permit persons to whom the Software
// is furnished to do so, subject to the following conditions:
// The above copyright notice and this permission notice shall be included in all copies or
// substantial portions of the Software.

////////////////////////////////////////////////////////////////////////////////
// Engineer:       Kerim TURAK - kerimturak@hotmail.com                       //
//                                                                            //
// Additional contributions by:                                               //
//                 --                                                         //
//                                                                            //
// Design Name:    dcache                                                     //
// Project Name:   TCORE                                                      //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    Writeback full configurable data cache                     //
////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
`include "tcore_defines.svh"
module dcache
  import tcore_param::*;
#(
    parameter CACHE_SIZE = (DC_CAPACITY),
    parameter BLK_SIZE = tcore_param::BLK_SIZE,
    parameter XLEN = tcore_param::XLEN,
    parameter NUM_WAY = DC_WAY
) (
    input  logic        clk_i,
    input  logic        rst_ni,
    input  dcache_req_t cache_req_i,
    output dcache_res_t cache_res_o,
    output logic        dcache_miss_o,
    input  dlowX_res_t  lowX_res_i,
    output dlowX_req_t  lowX_req_o
);

  localparam NUM_SET = (CACHE_SIZE / BLK_SIZE) / NUM_WAY;
  localparam IDX_WIDTH = $clog2(NUM_SET) == 0 ? 1 : $clog2(NUM_SET);
  localparam BOFFSET = $clog2(BLK_SIZE / 8);
  localparam WOFFSET = $clog2((BLK_SIZE / 32));
  localparam TAG_SIZE = XLEN - IDX_WIDTH - BOFFSET;

  logic                  cache_miss;
  logic                  cache_hit;
  logic  [IDX_WIDTH-1:0] pc_idx;
  logic  [  NUM_WAY-1:0] cache_wr_way;
  logic  [ BLK_SIZE-1:0] cache_select_data;
  logic  [ BLK_SIZE-1:0] mask_data;
  logic                  data_array_wr_en;
  logic  [ BLK_SIZE-1:0] data_wr_pre;
  logic  [ BLK_SIZE-1:0] data_wr_line;
  logic  [ BLK_SIZE-1:0] data_rd_line      [NUM_WAY];
  logic  [  NUM_WAY-1:0] data_write_way;
  logic                  tag_array_wr_en;
  logic  [   TAG_SIZE:0] cache_wr_tag;
  logic  [   TAG_SIZE:0] cache_rd_tag      [NUM_WAY];
  logic  [  NUM_WAY-1:0] evict_way;
  logic  [  NUM_WAY-1:0] cache_valid_vec;
  logic  [  NUM_WAY-1:0] cache_hit_vec;
  logic                  flush;
  logic  [IDX_WIDTH-1:0] flush_index;
  logic  [IDX_WIDTH-1:0] cache_idx;
  logic  [  NUM_WAY-1:0] tag_write_way;
  logic                  node_wr_en;
  logic  [  NUM_WAY-2:0] updated_node;
  logic  [  NUM_WAY-2:0] cache_wr_node;
  logic  [  NUM_WAY-2:0] cache_rd_node;
  logic  [  WOFFSET-1:0] word_idx;
  logic                  write_back;
  logic                  dirty_wr_en;
  logic  [  NUM_WAY-1:0] dirty_write_way;
  logic                  dirty_wr_data;
  logic  [  NUM_WAY-1:0] dirty_rd_data;
  logic  [ TAG_SIZE-1:0] evict_tag;
  logic  [ BLK_SIZE-1:0] evict_data;

  for (genvar i = 0; i < NUM_WAY; i++) begin : ddata_array
    sp_bram #(
        .DATA_WIDTH(BLK_SIZE),
        .NUM_SETS  (NUM_SET)
    ) data_array (
        .clk    (clk_i),
        .chip_en(1'b1),
        .addr   (pc_idx),
        .wr_en  (data_write_way[i]),
        .wr_data(data_wr_line),
        .rd_data(data_rd_line[i])
    );
  end

  for (genvar i = 0; i < NUM_WAY; i++) begin : dtag_array
    sp_bram #(
        .DATA_WIDTH(TAG_SIZE + 1),
        .NUM_SETS  (NUM_SET)
    ) tag_array (
        .clk    (clk_i),
        .chip_en(1'b1),
        .addr   (cache_idx),
        .wr_en  (tag_write_way[i]),
        .wr_data(cache_wr_tag),
        .rd_data(cache_rd_tag[i])
    );
  end

  for (genvar i = 0; i < NUM_WAY; i++) begin : ddirty_array
    sp_bram #(
        .DATA_WIDTH(1),
        .NUM_SETS  (NUM_SET)
    ) dirty_array (
        .clk    (clk_i),
        .chip_en(1'b1),
        .addr   (cache_idx),
        .wr_en  (dirty_write_way[i]),
        .wr_data(dirty_wr_data),
        .rd_data(dirty_rd_data[i])
    );
  end

  sp_bram #(
      .DATA_WIDTH(NUM_WAY - 1),
      .NUM_SETS  (NUM_SET)
  ) node_array (
      .clk    (clk_i),
      .chip_en(1'b1),
      .addr   (cache_idx),
      .wr_en  (node_wr_en),
      .wr_data(cache_wr_node),
      .rd_data(cache_rd_node)
  );

  plru #(
      .NUM_WAY(NUM_WAY)
  ) dplru (
      .node_i     (cache_rd_node),
      .hit_vec_i  (cache_hit_vec),
      .evict_way_o(evict_way),
      .node_o     (updated_node)
  );

  dcache_req_t cache_req_q;

  always_ff @(posedge clk_i) begin
    if (!rst_ni) begin
      cache_req_q <= '0;
      flush_index <= '0;
      flush       <= '1;
    end else begin
      cache_req_q      <= cache_req_i;
      if (flush && flush_index != 2 ** IDX_WIDTH - 1) begin
        flush_index <= flush_index + 1'b1;
      end else begin
        flush_index <= 1'b0;
        flush       <= 1'b0;
      end
    end
  end

  always_comb begin
    for (int i = 0; i < NUM_WAY; i++) begin
      cache_valid_vec[i] = cache_rd_tag[i][TAG_SIZE];
      cache_hit_vec[i]   = cache_rd_tag[i][TAG_SIZE-1:0] == cache_req_q.addr[XLEN-1:IDX_WIDTH+BOFFSET];
    end
    cache_wr_tag = flush ? '0 : {1'b1, cache_req_q.addr[XLEN-1:IDX_WIDTH+BOFFSET]};
    cache_wr_node = flush ? '0 : updated_node;
    cache_select_data = '0;
    for (int i = 0; i < NUM_WAY; i++) begin
      if (cache_hit_vec[i]) cache_select_data = data_rd_line[i];
    end
    cache_miss = cache_req_q.valid && !flush && !(|(cache_valid_vec & cache_hit_vec));
    cache_hit  = cache_req_q.valid && !flush &&  (|(cache_valid_vec & cache_hit_vec));

  end

  always_comb begin
    data_wr_pre = mask_data;
    case (cache_req_q.rw_size)
      WORD:      data_wr_pre[cache_req_i.addr[BOFFSET-1:2]*32+:32] = cache_req_q.data;
      HALF_WORD: data_wr_pre[cache_req_i.addr[BOFFSET-1:1]*16+:16] = cache_req_q.data;
      BYTE:      data_wr_pre[cache_req_i.addr[BOFFSET-1:0]*8+:8] = cache_req_q.data;
      NO_SIZE:   data_wr_pre = '0;
    endcase
  end

  always_comb begin
    write_back = cache_miss && (|(dirty_rd_data & evict_way & cache_valid_vec));


    data_array_wr_en = (cache_hit && cache_req_q.rw) || (cache_miss && lowX_res_i.valid && !cache_req_q.uncached) && !write_back; // icachte cache_wr_En'e denk
    tag_array_wr_en = (cache_miss && lowX_res_i.valid && !cache_req_q.uncached) && !write_back;
    node_wr_en    = flush || data_array_wr_en;
    cache_wr_way = cache_hit ? cache_hit_vec : evict_way;


    for (int i = 0; i < NUM_WAY; i++) data_write_way[i] = cache_wr_way[i] && data_array_wr_en;
    for (int i = 0; i < NUM_WAY; i++) tag_write_way[i] = flush ? '1 : cache_wr_way[i] && tag_array_wr_en || flush;



    pc_idx = cache_req_i.addr[IDX_WIDTH+BOFFSET:BOFFSET];
    cache_idx = flush ? flush_index : pc_idx;

    dirty_wr_en = (cache_req_q.rw && (cache_hit || (cache_miss && lowX_res_i.valid))) || (write_back && lowX_res_i.valid);
    for (int i = 0; i < NUM_WAY; i++) dirty_write_way[i] = flush ? '1 : cache_wr_way[i] && dirty_wr_en || flush;
    dirty_wr_data = flush ? '0 : (write_back ? '0 : cache_req_q.rw ? '1 : '0);

    evict_tag = '0;
    evict_data = '0;
    for (int i = 0; i < NUM_WAY; i++) if (evict_way[i]) evict_tag = cache_rd_tag[i][TAG_SIZE-1:0];
    for (int i = 0; i < NUM_WAY; i++) if (evict_way[i]) evict_data = data_rd_line[i];


    mask_data = cache_hit ? cache_select_data : lowX_res_i.data;
    data_wr_line = cache_req_q.rw ? data_wr_pre : lowX_res_i.data;

  end

  always_comb begin
    word_idx = cache_req_i.addr[(WOFFSET+2)-1:2];
    lowX_req_o.valid = cache_miss && lowX_res_i.ready;
    lowX_req_o.ready = 1'b1;
    lowX_req_o.uncached = write_back ? '0 : cache_req_q.uncached;
    lowX_req_o.addr = write_back ? {evict_tag, pc_idx, {BOFFSET{1'b0}}} : {cache_req_q.addr[31:BOFFSET], {BOFFSET{1'b0}}};
    lowX_req_o.rw = write_back ? '1 : '0;
    lowX_req_o.rw_size = write_back ? WORD : cache_req_q.rw_size;
    lowX_req_o.data = write_back ? evict_data : '0;

    cache_res_o.valid = !cache_req_q.rw ? !write_back && cache_req_q.valid &&  (cache_hit || (cache_miss && lowX_req_o.ready && lowX_res_i.valid)) :
                        !write_back && cache_req_q.valid && cache_req_i.ready  && (cache_hit || (cache_miss && lowX_req_o.ready && lowX_res_i.valid));
    cache_res_o.ready = !cache_req_q.rw ? !write_back && (!cache_miss || lowX_res_i.valid) && !flush && !tag_array_wr_en : !write_back && !tag_array_wr_en && lowX_req_o.ready && lowX_res_i.valid && !flush;
    dcache_miss_o = cache_miss;
    cache_res_o.data = (cache_miss && lowX_res_i.valid) ? lowX_res_i.data[word_idx*32+:32] : cache_select_data[word_idx*32+:32];
  end

endmodule
