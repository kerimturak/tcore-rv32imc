//`define STATIC_PREDICT
`define RAS
//`define WALLACE_SINGLE_CYCLE
//`define WALLACE_MULTY_CYCLE
`define DSP_MUL
//`define REMOVE_WB_STAGE