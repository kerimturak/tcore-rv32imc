package configure;
  timeunit 1ps;
  timeprecision 1ps;

  parameter XLEN = 32;
  parameter YLEN = 32;
  parameter TYP = 0;
  integer MAXTIME = 10;
  integer SEED = 1722709091;
endpackage
